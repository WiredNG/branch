`ifndef _BRPACKAGES
`define _BRPACKAGES
import WiredSpec::*;
import WiredL1BTB::*;
import WiredTAGE::*;
import WiredBranchDefines::*;
`endif
